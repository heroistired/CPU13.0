library verilog;
use verilog.vl_types.all;
entity systemC is
    port(
        writemem        : out    vl_logic;
        flagin          : out    vl_logic_vector(1 downto 0);
        flagout         : out    vl_logic_vector(7 downto 0);
        CLK             : in     vl_logic;
        RST             : in     vl_logic;
        wrflag          : out    vl_logic;
        cs              : out    vl_logic_vector(3 downto 0);
        Q1              : out    vl_logic_vector(7 downto 0);
        reg_we          : out    vl_logic;
        DI              : out    vl_logic_vector(7 downto 0);
        memtoreg        : out    vl_logic;
        S               : out    vl_logic_vector(7 downto 0);
        ram             : out    vl_logic_vector(7 downto 0);
        io_read         : out    vl_logic;
        Q2              : out    vl_logic_vector(7 downto 0);
        V               : out    vl_logic_vector(3 downto 0);
        H               : out    vl_logic_vector(3 downto 0);
        key             : in     vl_logic_vector(15 downto 0);
        instr           : out    vl_logic_vector(15 downto 0);
        pc              : out    vl_logic_vector(7 downto 0);
        branch          : out    vl_logic;
        jump            : out    vl_logic;
        ND              : out    vl_logic_vector(7 downto 0);
        regdes          : out    vl_logic;
        ALUSRCB         : out    vl_logic;
        sign            : out    vl_logic;
        AALU_OP         : out    vl_logic_vector(7 downto 0);
        data_inH        : out    vl_logic_vector(7 downto 0);
        data_inL        : out    vl_logic_vector(7 downto 0);
        data_out        : out    vl_logic_vector(7 downto 0);
        DSTH            : out    vl_logic_vector(7 downto 0);
        DSTL            : out    vl_logic_vector(7 downto 0);
        finish_sign     : out    vl_logic_vector(7 downto 0);
        IO0             : out    vl_logic_vector(7 downto 0);
        IO1             : out    vl_logic_vector(7 downto 0);
        N1              : out    vl_logic_vector(1 downto 0);
        N2              : out    vl_logic_vector(1 downto 0);
        num_C0          : out    vl_logic_vector(3 downto 0);
        num_C1          : out    vl_logic_vector(3 downto 0);
        num_C2          : out    vl_logic_vector(3 downto 0);
        num_C3          : out    vl_logic_vector(3 downto 0);
        result          : out    vl_logic_vector(7 downto 0);
        seg_sel         : out    vl_logic_vector(3 downto 0);
        SRCH            : out    vl_logic_vector(7 downto 0);
        SRCL            : out    vl_logic_vector(7 downto 0)
    );
end systemC;
