library verilog;
use verilog.vl_types.all;
entity IO_PORT_vlg_vec_tst is
end IO_PORT_vlg_vec_tst;
