library verilog;
use verilog.vl_types.all;
entity instrconunit_vlg_vec_tst is
end instrconunit_vlg_vec_tst;
