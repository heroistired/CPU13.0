library verilog;
use verilog.vl_types.all;
entity systemC_vlg_vec_tst is
end systemC_vlg_vec_tst;
