library verilog;
use verilog.vl_types.all;
entity alu8_vlg_vec_tst is
end alu8_vlg_vec_tst;
