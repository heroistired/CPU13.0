library verilog;
use verilog.vl_types.all;
entity ctrlunit_vlg_vec_tst is
end ctrlunit_vlg_vec_tst;
