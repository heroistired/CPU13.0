library verilog;
use verilog.vl_types.all;
entity NixieScan_vlg_vec_tst is
end NixieScan_vlg_vec_tst;
