library verilog;
use verilog.vl_types.all;
entity myrom_vlg_vec_tst is
end myrom_vlg_vec_tst;
