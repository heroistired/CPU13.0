library verilog;
use verilog.vl_types.all;
entity lpm_rom_256_16_vlg_vec_tst is
end lpm_rom_256_16_vlg_vec_tst;
