library verilog;
use verilog.vl_types.all;
entity myram_256_8_vlg_vec_tst is
end myram_256_8_vlg_vec_tst;
