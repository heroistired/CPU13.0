library verilog;
use verilog.vl_types.all;
entity systemB_vlg_vec_tst is
end systemB_vlg_vec_tst;
