library verilog;
use verilog.vl_types.all;
entity systemA_vlg_vec_tst is
end systemA_vlg_vec_tst;
