library verilog;
use verilog.vl_types.all;
entity systemB_vlg_check_tst is
    port(
        ALUSRCB         : in     vl_logic;
        branch          : in     vl_logic;
        cs              : in     vl_logic_vector(3 downto 0);
        data_inH        : in     vl_logic_vector(7 downto 0);
        data_inL        : in     vl_logic_vector(7 downto 0);
        DI              : in     vl_logic_vector(7 downto 0);
        flagin          : in     vl_logic_vector(1 downto 0);
        flagout         : in     vl_logic_vector(7 downto 0);
        instr           : in     vl_logic_vector(15 downto 0);
        IO0             : in     vl_logic_vector(7 downto 0);
        IO1             : in     vl_logic_vector(7 downto 0);
        IO_read         : in     vl_logic;
        jump            : in     vl_logic;
        memtoreg        : in     vl_logic;
        N1              : in     vl_logic_vector(1 downto 0);
        N2              : in     vl_logic_vector(1 downto 0);
        ND              : in     vl_logic_vector(7 downto 0);
        num_C0          : in     vl_logic_vector(3 downto 0);
        num_C1          : in     vl_logic_vector(3 downto 0);
        num_C2          : in     vl_logic_vector(3 downto 0);
        num_C3          : in     vl_logic_vector(3 downto 0);
        pc              : in     vl_logic_vector(7 downto 0);
        q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        q3              : in     vl_logic;
        q4              : in     vl_logic;
        q5              : in     vl_logic;
        q6              : in     vl_logic;
        q7              : in     vl_logic;
        Q10             : in     vl_logic;
        Q11             : in     vl_logic;
        Q12             : in     vl_logic;
        Q13             : in     vl_logic;
        Q14             : in     vl_logic;
        Q15             : in     vl_logic;
        Q16             : in     vl_logic;
        Q17             : in     vl_logic;
        Q20             : in     vl_logic;
        Q21             : in     vl_logic;
        Q22             : in     vl_logic;
        Q23             : in     vl_logic;
        Q24             : in     vl_logic;
        Q25             : in     vl_logic;
        Q26             : in     vl_logic;
        Q27             : in     vl_logic;
        ram             : in     vl_logic_vector(7 downto 0);
        reg_we          : in     vl_logic;
        regdes          : in     vl_logic;
        result          : in     vl_logic_vector(7 downto 0);
        S               : in     vl_logic_vector(7 downto 0);
        sign            : in     vl_logic;
        wrflag          : in     vl_logic;
        writemem        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end systemB_vlg_check_tst;
